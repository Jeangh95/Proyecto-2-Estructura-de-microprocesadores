`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.08.2017 08:51:36
// Design Name: 
// Module Name: Mux_EN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mux_EN(out_mux,sel_mux);
output reg [31:0]out_mux;
input  [0:4]sel_mux;

always @ (sel_mux or out_mux)
case(sel_mux)
5'b00000: out_mux=32'b00000000000000000000000000000001;
5'b00001: out_mux=32'b00000000000000000000000000000010;
5'b00010: out_mux=32'b00000000000000000000000000000100;
5'b00011: out_mux=32'b00000000000000000000000000001000;
5'b00100: out_mux=32'b00000000000000000000000000010000;
5'b00101: out_mux=32'b00000000000000000000000000100000;
5'b00110: out_mux=32'b00000000000000000000000001000000;
5'b00111: out_mux=32'b00000000000000000000000010000000;
5'b01000: out_mux=32'b00000000000000000000000100000000;
5'b01001: out_mux=32'b00000000000000000000001000000000;
5'b01010: out_mux=32'b00000000000000000000010000000000;
5'b01011: out_mux=32'b00000000000000000000100000000000;
5'b01100: out_mux=32'b00000000000000000001000000000000;
5'b01101: out_mux=32'b00000000000000000010000000000000;
5'b01110: out_mux=32'b00000000000000000100000000000000;
5'b01111: out_mux=32'b00000000000000001000000000000000;
5'b10000: out_mux=32'b00000000000000010000000000000000;
5'b10001: out_mux=32'b00000000000000100000000000000000;
5'b10010: out_mux=32'b00000000000001000000000000000000;
5'b10011: out_mux=32'b00000000000010000000000000000000;
5'b10100: out_mux=32'b00000000000100000000000000000000;
5'b10101: out_mux=32'b00000000001000000000000000000000;
5'b10110: out_mux=32'b00000000010000000000000000000000;
5'b10111: out_mux=32'b00000000100000000000000000000000;
5'b11000: out_mux=32'b00000001000000000000000000000000;
5'b11001: out_mux=32'b00000010000000000000000000000000;
5'b11010: out_mux=32'b00000100000000000000000000000000;
5'b11011: out_mux=32'b00001000000000000000000000000000;
5'b11100: out_mux=32'b00010000000000000000000000000000;
5'b11101: out_mux=32'b00100000000000000000000000000000;
5'b11110: out_mux=32'b01000000000000000000000000000000;
5'b11111: out_mux=32'b10000000000000000000000000000000;
endcase
endmodule